-------------------------------------------------------------------------------
-- Title      : LoRa core
-- Project    : Travail de bachelor
-------------------------------------------------------------------------------
-- File       : lora_detect.vhd
-- Author     :   <seba@t440p>
-- Company    : HESSO - hepia - ITI
-- Created    : 2017-06-18
-- Last update: 2017-06-20
-- Platform   :
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: This module detect a LoRa packet in a stream of data from an
--              ADC and timestamp it.
-------------------------------------------------------------------------------
-- Copyright (c) 2017 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2017-05-17  1.0      seba  Created
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity lora_detect is

--    generic (
--        NB_OF_SAMPLES : 64);            -- sample

  port (
    -- TODO choose one clock
    radio_clk : in std_logic;           -- radio clock 
    bus_clk   : in std_logic;           -- bus clock
    rst       : in std_logic;           -- reset SR registers

    rx_i      : in std_logic_vector(15 downto 0);  -- rx I signal
    rx_q      : in std_logic_vector(15 downto 0);  -- rx Q signal
    vita_time : in std_logic_vector(63 downto 0);  -- vita time
    trigger_i : in std_logic;                      -- external trigger

    -- wishbone
    addr   : in std_logic_vector(7 downto 0);   -- setting reg
    data   : in std_logic_vector(31 downto 0);  -- data
    strobe : in std_logic;

    -- debug chipscope
    chipscope_bus_o     : out std_logic_vector(5 downto 0);  -- probe chipscope
    chipscope_radio_o   : out std_logic_vector(33 downto 0);  -- probe chipscope
    -- readback output
    lora_time_measured_o : out std_logic_vector(63 downto 0));  -- detected packet's trigger

end entity lora_detect;

architecture lora_detect_behav of lora_detect is

  ------------------------------------
  -- Components
  ------------------------------------
  component gen_event_trigger is
    port (
      clk       : in std_logic;
      rst       : in std_logic;
      trigger_i : in std_logic);
  end component gen_event_trigger;

  component setting_reg_vhdl_wrapper is
    port (
      clk      : in  std_logic;
      rst      : in  std_logic;
      strobe   : in  std_logic;
      addr     : in  std_logic_vector(7 downto 0);
      data_in  : in  std_logic_vector(31 downto 0);
      data_out : out std_logic_vector(31 downto 0));
  end component setting_reg_vhdl_wrapper;


  -------------------------------------------------------
  -- signals
  -------------------------------------------------------
  signal sr0_value_int     : std_logic_vector(31 downto 0);  -- setting register value
  signal sr0_value_nxt_int : std_logic_vector(31 downto 0);  -- setting register value

  signal save_time_int        : std_logic := '0';  -- enable measure
  signal gen_soft_trigger_int : std_logic;         -- lora detected
  signal gen_uart_trigger_int : std_logic;         -- trigger rising edge
  signal gen_lora_trigger_int : std_logic := '0';  -- trigger rising edge


begin  -- architecture lora_detect_behav

  --------------------------
  -- setting register 0
  -- cpp API trigger
  --------------------------
  sr_lora_0 : setting_reg_vhdl_wrapper port map (
    clk      => bus_clk,
    rst      => rst,
    strobe   => strobe,
    addr     => addr,
    data_in  => data,
    data_out => sr0_value_int);

  --------------------------------
  -- Enable register vita time
  -- combinational
  --------------------------------
  save_time_int <= gen_lora_trigger_int or gen_soft_trigger_int or gen_uart_trigger_int;

  -----------------------------------
  -- instance "gen_event_trigger_1"
  -----------------------------------
  gen_uart_trigger_1 : entity work.gen_event_trigger
    port map (
      clk       => radio_clk,
      rst       => rst,
      trigger_i => trigger_i,
      trigger_o => gen_uart_trigger_int);

  -----------------------------------
  -- instance "gen_soft_trigger_1"
  -----------------------------------
  gen_soft_trigger_1 : entity work.gen_event_trigger
    port map (
      clk       => bus_clk,
      rst       => rst,
      trigger_i => sr0_value_int(0),
      trigger_o => gen_soft_trigger_int);

  -----------------------------------
  -- instance "gen_lora_trigger_1"
  -----------------------------------
  -- gen_lora_trigger_1 : entity work.gen_event_trigger
  --   port map (
  --     clk       => bus_clk,
  --     rst       => rst,
  --     trigger_i => lora_i,
  --     trigger_o => gen_lora_trigger_int);

  ----------------------------------------
  -- purpose: one cycle only trigger
  -- type   : sequential
  -- inputs : bus_clk, rst, sr0_value_int
  -- outputs: one pulse when register ==0x1
  ----------------------------------------
  -- software_trig : process (bus_clk, rst) is
  -- begin  -- process measure
  --   if rst = '1' then                   -- asynchronous reset (active low)
  --   --sr0_value_int <= (others => '0');
  --   elsif rising_edge(bus_clk) then     -- rising clock edge
  --     sr0_value_nxt_int <= sr0_value_int;
  --   end if;
  -- end process software_trig;

  -- gen_soft_trigger_int <= '1' when sr0_value_nxt_int(0) = '0' and sr0_value_int(0) = '1' else '0';

----------------------------------------
-- purpose: timestamp register
-- type   : sequential
-- inputs : bus_clk, rst, en_measure_int
-- outputs: measured_time
----------------------------------------
  measure : process (radio_clk, rst) is
  begin  -- process measure
    if rst = '0' then                   -- asynchronous reset (active low)
      lora_time_measured_o <= (others => '0');
    elsif rising_edge(radio_clk) then   -- rising clock edge
      if save_time_int = '1' then
        lora_time_measured_o <= vita_time;
      end if;
    end if;
  end process measure;

--------------------------------------
-- Debug with chipscope
--------------------------------------
  --chipscope_o <= ( rx_q & rx_i & "000000000" & strobe & rst & save_time_int & gen_lora_trigger_int & gen_soft_trigger_int & gen_uart_trigger_int & trigger_i & sr0_value_int(7 downto 0) & addr);
  chipscope_bus_o <= ('0' & strobe & rst & save_time_int & gen_lora_trigger_int & gen_soft_trigger_int);
  chipscope_radio_o <= (rx_q & rx_i & gen_uart_trigger_int & trigger_i);

-- 4 pps avant et aprs mux            (4bits)
-- strobe, rst, soft_trig, save, uart  (4bits)
-- rx i/q                             (32bits)
-- rb_data et set_data[7:0]           (16bits)
-- set_addr et rb_addr                (16bits)
-- vita[31:0] et vita_reg[31:0]       (64bits)
-- 
end architecture lora_detect_behav;
