seba@t440p.4053:1497801611